liBRARy ieee; uSE Ieee.STd_LOgIC_1164.ALL; eNtIty iD_S_b88a693_7e3412F0_e iS pORt( iD_S_B88665F_7e7082e6_e : In Std_logiC; Id_S_59777b_7FFCe7eC_E : In sTD_LoGIc; id_s_c89sdnc7u_sda09scah_E : iN STd_lOGic; id_s_daf34r31df1d_0y8wefh80_E : iN STd_Logic_vECtoR(9 DoWNto 0); ID_S_191530b5_24e2B0Bf_E : OuT sTd_LOGIc_vECtoR(31 DowNTo 0) ); End iD_s_B88A693_7E3412f0_e; ARchITectURe id_s_455b727d_1f58D85f_e of id_s_B88a693_7E3412f0_E Is cOMPonent ROM_Block is pORT( address : In sTd_LOGIC_vEctOR(9 DoWnTO 0); clOCK : In sTD_loGIc; q : oUT sTD_LoGic_VeCTor(31 downTO 0) ); EnD ComponeNT; SigNAL Id_s_515D507a_5d491c3b_E : std_LOGic_veCTOR(31 dOWNTO 0); siGNAl Id_S_294e5c0d_762308e6_E : std_loGIc; BeGIN iD_s_30739CAe_5A20DAf5_E : ROM_Block porT mAp( address => id_s_daf34r31df1d_0y8wefh80_E, CLOck => id_s_b88665F_7e7082e6_E, q => ID_s_515D507A_5d491C3b_E ); PROCESs(id_s_B88665f_7e7082E6_e) beGIN If (risiNg_EDGE(id_S_b88665F_7e7082E6_e)) TheN ID_s_294e5c0D_762308E6_E <= id_s_c89sdnc7u_sda09scah_E and iD_S_59777B_7fFCE7EC_E; eNd iF; ENd pROceSS; PrOCESS(id_S_294e5C0d_762308E6_E, id_S_515d507a_5d491C3b_E) bEgiN Id_S_191530B5_24E2b0Bf_E <= (others => 'Z'); iF ( ID_s_294E5c0D_762308e6_E = '1') THeN ID_S_191530B5_24e2b0BF_E <= iD_s_515D507a_5D491C3b_E; EnD IF; End proceSS; eNd iD_s_455B727D_1f58D85f_e;